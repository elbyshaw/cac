module tb_systolic;
	parameter CLK_PERIOD = 10;


endmodule

