package pkg;
    parameter NUM_BITS = 8;

    typedef enum logic [1:0] {S_PASSTHROUGH,S_LOAD,S_PROCESS} input_mux_t;
    //TODO: Add any typedefs, enums, or parameters as neccessary for your project

endpackage