
module
	input top
	input left
	
	output right
	output bottom

endmodule
